** sch_path: /pri/bjs1/aicex/ip/jnw_bkle_sky130A/design/JNW_BKLE_SKY130A/JNW_BKLE.sch
**.subckt JNW_BKLE IBPS_2U VSS IBNS_20U
*.ipin IBPS_2U
*.ipin VSS
*.ipin IBNS_20U
x1 IBNS_20U IBPS_2U VSS VSS JNWATR_NCH_12C1F2
x2 IBPS_2U IBPS_2U VSS VSS JNWATR_NCH_2C1F2
**.ends

* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_12C1F2.sym # of pins=4
** sym_path: /pri/bjs1/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A/JNWATR_NCH_12C1F2.sym
** sch_path: /pri/bjs1/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A/JNWATR_NCH_12C1F2.sch
.subckt JNWATR_NCH_12C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=8.32 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym # of pins=4
** sym_path: /pri/bjs1/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym
** sch_path: /pri/bjs1/aicex/ip/jnw_bkle_sky130A/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sch
.subckt JNWATR_NCH_2C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=1.92 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
